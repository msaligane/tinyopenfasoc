magic
tech sky130A
magscale 1 2
timestamp 1662472490
<< viali >>
rect 25421 47141 25455 47175
rect 1409 47073 1443 47107
rect 1685 47005 1719 47039
rect 25237 47005 25271 47039
rect 48053 37825 48087 37859
rect 47961 37621 47995 37655
rect 24501 25857 24535 25891
rect 25053 25857 25087 25891
rect 24961 25789 24995 25823
rect 24317 25653 24351 25687
rect 41337 25449 41371 25483
rect 41521 25245 41555 25279
rect 48145 25245 48179 25279
rect 47961 25109 47995 25143
rect 41521 24837 41555 24871
rect 1593 24769 1627 24803
rect 2237 24769 2271 24803
rect 25053 24769 25087 24803
rect 25513 24769 25547 24803
rect 41797 24769 41831 24803
rect 47869 24769 47903 24803
rect 2421 24633 2455 24667
rect 24869 24633 24903 24667
rect 48053 24633 48087 24667
rect 1777 24565 1811 24599
rect 25697 24565 25731 24599
rect 47869 24361 47903 24395
rect 1777 24157 1811 24191
rect 47869 24157 47903 24191
rect 1593 24021 1627 24055
rect 24869 7837 24903 7871
rect 25053 7701 25087 7735
rect 1593 2601 1627 2635
rect 37565 2465 37599 2499
rect 46765 2465 46799 2499
rect 1409 2397 1443 2431
rect 12357 2397 12391 2431
rect 37289 2397 37323 2431
rect 47041 2397 47075 2431
rect 12541 2261 12575 2295
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 25409 47175 25467 47181
rect 25409 47141 25421 47175
rect 25455 47172 25467 47175
rect 25498 47172 25504 47184
rect 25455 47144 25504 47172
rect 25455 47141 25467 47144
rect 25409 47135 25467 47141
rect 25498 47132 25504 47144
rect 25556 47132 25562 47184
rect 658 47064 664 47116
rect 716 47104 722 47116
rect 1397 47107 1455 47113
rect 1397 47104 1409 47107
rect 716 47076 1409 47104
rect 716 47064 722 47076
rect 1397 47073 1409 47076
rect 1443 47073 1455 47107
rect 1397 47067 1455 47073
rect 1578 46996 1584 47048
rect 1636 47036 1642 47048
rect 1673 47039 1731 47045
rect 1673 47036 1685 47039
rect 1636 47008 1685 47036
rect 1636 46996 1642 47008
rect 1673 47005 1685 47008
rect 1719 47005 1731 47039
rect 25222 47036 25228 47048
rect 25183 47008 25228 47036
rect 1673 46999 1731 47005
rect 25222 46996 25228 47008
rect 25280 46996 25286 47048
rect 37366 46860 37372 46912
rect 37424 46900 37430 46912
rect 39298 46900 39304 46912
rect 37424 46872 39304 46900
rect 37424 46860 37430 46872
rect 39298 46860 39304 46872
rect 39356 46860 39362 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 48130 46044 48136 46096
rect 48188 46084 48194 46096
rect 49602 46084 49608 46096
rect 48188 46056 49608 46084
rect 48188 46044 48194 46056
rect 49602 46044 49608 46056
rect 49660 46044 49666 46096
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 48038 37856 48044 37868
rect 47999 37828 48044 37856
rect 48038 37816 48044 37828
rect 48096 37816 48102 37868
rect 25038 37612 25044 37664
rect 25096 37652 25102 37664
rect 47949 37655 48007 37661
rect 47949 37652 47961 37655
rect 25096 37624 47961 37652
rect 25096 37612 25102 37624
rect 47949 37621 47961 37624
rect 47995 37621 48007 37655
rect 47949 37615 48007 37621
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 24489 25891 24547 25897
rect 24489 25857 24501 25891
rect 24535 25857 24547 25891
rect 25038 25888 25044 25900
rect 24999 25860 25044 25888
rect 24489 25851 24547 25857
rect 24504 25820 24532 25851
rect 25038 25848 25044 25860
rect 25096 25848 25102 25900
rect 24949 25823 25007 25829
rect 24949 25820 24961 25823
rect 24504 25792 24961 25820
rect 24949 25789 24961 25792
rect 24995 25789 25007 25823
rect 24949 25783 25007 25789
rect 3418 25644 3424 25696
rect 3476 25684 3482 25696
rect 24305 25687 24363 25693
rect 24305 25684 24317 25687
rect 3476 25656 24317 25684
rect 3476 25644 3482 25656
rect 24305 25653 24317 25656
rect 24351 25653 24363 25687
rect 24305 25647 24363 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 39298 25440 39304 25492
rect 39356 25480 39362 25492
rect 41325 25483 41383 25489
rect 41325 25480 41337 25483
rect 39356 25452 41337 25480
rect 39356 25440 39362 25452
rect 41325 25449 41337 25452
rect 41371 25449 41383 25483
rect 41325 25443 41383 25449
rect 41506 25276 41512 25288
rect 41467 25248 41512 25276
rect 41506 25236 41512 25248
rect 41564 25236 41570 25288
rect 48130 25276 48136 25288
rect 48091 25248 48136 25276
rect 48130 25236 48136 25248
rect 48188 25236 48194 25288
rect 46750 25100 46756 25152
rect 46808 25140 46814 25152
rect 47949 25143 48007 25149
rect 47949 25140 47961 25143
rect 46808 25112 47961 25140
rect 46808 25100 46814 25112
rect 47949 25109 47961 25112
rect 47995 25109 48007 25143
rect 47949 25103 48007 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 41506 24868 41512 24880
rect 41467 24840 41512 24868
rect 41506 24828 41512 24840
rect 41564 24828 41570 24880
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 2225 24803 2283 24809
rect 2225 24769 2237 24803
rect 2271 24769 2283 24803
rect 25038 24800 25044 24812
rect 24999 24772 25044 24800
rect 2225 24763 2283 24769
rect 1486 24692 1492 24744
rect 1544 24732 1550 24744
rect 2240 24732 2268 24763
rect 25038 24760 25044 24772
rect 25096 24760 25102 24812
rect 25498 24800 25504 24812
rect 25459 24772 25504 24800
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 41785 24803 41843 24809
rect 41785 24769 41797 24803
rect 41831 24800 41843 24803
rect 46750 24800 46756 24812
rect 41831 24772 46756 24800
rect 41831 24769 41843 24772
rect 41785 24763 41843 24769
rect 46750 24760 46756 24772
rect 46808 24760 46814 24812
rect 47854 24800 47860 24812
rect 47815 24772 47860 24800
rect 47854 24760 47860 24772
rect 47912 24760 47918 24812
rect 1544 24704 2268 24732
rect 1544 24692 1550 24704
rect 2406 24664 2412 24676
rect 2367 24636 2412 24664
rect 2406 24624 2412 24636
rect 2464 24624 2470 24676
rect 12434 24624 12440 24676
rect 12492 24664 12498 24676
rect 24857 24667 24915 24673
rect 24857 24664 24869 24667
rect 12492 24636 24869 24664
rect 12492 24624 12498 24636
rect 24857 24633 24869 24636
rect 24903 24633 24915 24667
rect 48038 24664 48044 24676
rect 47999 24636 48044 24664
rect 24857 24627 24915 24633
rect 48038 24624 48044 24636
rect 48096 24624 48102 24676
rect 1762 24596 1768 24608
rect 1723 24568 1768 24596
rect 1762 24556 1768 24568
rect 1820 24556 1826 24608
rect 23474 24556 23480 24608
rect 23532 24596 23538 24608
rect 25685 24599 25743 24605
rect 25685 24596 25697 24599
rect 23532 24568 25697 24596
rect 23532 24556 23538 24568
rect 25685 24565 25697 24568
rect 25731 24565 25743 24599
rect 25685 24559 25743 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 47854 24392 47860 24404
rect 47815 24364 47860 24392
rect 47854 24352 47860 24364
rect 47912 24352 47918 24404
rect 1762 24188 1768 24200
rect 1723 24160 1768 24188
rect 1762 24148 1768 24160
rect 1820 24148 1826 24200
rect 47854 24188 47860 24200
rect 47815 24160 47860 24188
rect 47854 24148 47860 24160
rect 47912 24148 47918 24200
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24052 1639 24055
rect 2774 24052 2780 24064
rect 1627 24024 2780 24052
rect 1627 24021 1639 24024
rect 1581 24015 1639 24021
rect 2774 24012 2780 24024
rect 2832 24012 2838 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 20254 7828 20260 7880
rect 20312 7868 20318 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 20312 7840 24869 7868
rect 20312 7828 20318 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 25041 7735 25099 7741
rect 25041 7701 25053 7735
rect 25087 7732 25099 7735
rect 46382 7732 46388 7744
rect 25087 7704 46388 7732
rect 25087 7701 25099 7704
rect 25041 7695 25099 7701
rect 46382 7692 46388 7704
rect 46440 7692 46446 7744
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 1486 2592 1492 2644
rect 1544 2632 1550 2644
rect 1581 2635 1639 2641
rect 1581 2632 1593 2635
rect 1544 2604 1593 2632
rect 1544 2592 1550 2604
rect 1581 2601 1593 2604
rect 1627 2601 1639 2635
rect 1581 2595 1639 2601
rect 37553 2499 37611 2505
rect 37553 2496 37565 2499
rect 26206 2468 37565 2496
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12308 2400 12357 2428
rect 12308 2388 12314 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 25038 2388 25044 2440
rect 25096 2428 25102 2440
rect 26206 2428 26234 2468
rect 37553 2465 37565 2468
rect 37599 2465 37611 2499
rect 37553 2459 37611 2465
rect 46753 2499 46811 2505
rect 46753 2465 46765 2499
rect 46799 2496 46811 2499
rect 47854 2496 47860 2508
rect 46799 2468 47860 2496
rect 46799 2465 46811 2468
rect 46753 2459 46811 2465
rect 47854 2456 47860 2468
rect 47912 2456 47918 2508
rect 25096 2400 26234 2428
rect 25096 2388 25102 2400
rect 36722 2388 36728 2440
rect 36780 2428 36786 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36780 2400 37289 2428
rect 36780 2388 36786 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 47029 2431 47087 2437
rect 47029 2397 47041 2431
rect 47075 2428 47087 2431
rect 48958 2428 48964 2440
rect 47075 2400 48964 2428
rect 47075 2397 47087 2400
rect 47029 2391 47087 2397
rect 48958 2388 48964 2400
rect 49016 2388 49022 2440
rect 12529 2295 12587 2301
rect 12529 2261 12541 2295
rect 12575 2292 12587 2295
rect 20254 2292 20260 2304
rect 12575 2264 20260 2292
rect 12575 2261 12587 2264
rect 12529 2255 12587 2261
rect 20254 2252 20260 2264
rect 20312 2252 20318 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 25504 47132 25556 47184
rect 664 47064 716 47116
rect 1584 46996 1636 47048
rect 25228 47039 25280 47048
rect 25228 47005 25237 47039
rect 25237 47005 25271 47039
rect 25271 47005 25280 47039
rect 25228 46996 25280 47005
rect 37372 46860 37424 46912
rect 39304 46860 39356 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 48136 46044 48188 46096
rect 49608 46044 49660 46096
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 48044 37859 48096 37868
rect 48044 37825 48053 37859
rect 48053 37825 48087 37859
rect 48087 37825 48096 37859
rect 48044 37816 48096 37825
rect 25044 37612 25096 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 25044 25891 25096 25900
rect 25044 25857 25053 25891
rect 25053 25857 25087 25891
rect 25087 25857 25096 25891
rect 25044 25848 25096 25857
rect 3424 25644 3476 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 39304 25440 39356 25492
rect 41512 25279 41564 25288
rect 41512 25245 41521 25279
rect 41521 25245 41555 25279
rect 41555 25245 41564 25279
rect 41512 25236 41564 25245
rect 48136 25279 48188 25288
rect 48136 25245 48145 25279
rect 48145 25245 48179 25279
rect 48179 25245 48188 25279
rect 48136 25236 48188 25245
rect 46756 25100 46808 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 41512 24871 41564 24880
rect 41512 24837 41521 24871
rect 41521 24837 41555 24871
rect 41555 24837 41564 24871
rect 41512 24828 41564 24837
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 25044 24803 25096 24812
rect 1492 24692 1544 24744
rect 25044 24769 25053 24803
rect 25053 24769 25087 24803
rect 25087 24769 25096 24803
rect 25044 24760 25096 24769
rect 25504 24803 25556 24812
rect 25504 24769 25513 24803
rect 25513 24769 25547 24803
rect 25547 24769 25556 24803
rect 25504 24760 25556 24769
rect 46756 24760 46808 24812
rect 47860 24803 47912 24812
rect 47860 24769 47869 24803
rect 47869 24769 47903 24803
rect 47903 24769 47912 24803
rect 47860 24760 47912 24769
rect 2412 24667 2464 24676
rect 2412 24633 2421 24667
rect 2421 24633 2455 24667
rect 2455 24633 2464 24667
rect 2412 24624 2464 24633
rect 12440 24624 12492 24676
rect 48044 24667 48096 24676
rect 48044 24633 48053 24667
rect 48053 24633 48087 24667
rect 48087 24633 48096 24667
rect 48044 24624 48096 24633
rect 1768 24599 1820 24608
rect 1768 24565 1777 24599
rect 1777 24565 1811 24599
rect 1811 24565 1820 24599
rect 1768 24556 1820 24565
rect 23480 24556 23532 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 47860 24395 47912 24404
rect 47860 24361 47869 24395
rect 47869 24361 47903 24395
rect 47903 24361 47912 24395
rect 47860 24352 47912 24361
rect 1768 24191 1820 24200
rect 1768 24157 1777 24191
rect 1777 24157 1811 24191
rect 1811 24157 1820 24191
rect 1768 24148 1820 24157
rect 47860 24191 47912 24200
rect 47860 24157 47869 24191
rect 47869 24157 47903 24191
rect 47903 24157 47912 24191
rect 47860 24148 47912 24157
rect 2780 24012 2832 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 20260 7828 20312 7880
rect 46388 7692 46440 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1492 2592 1544 2644
rect 20 2388 72 2440
rect 12256 2388 12308 2440
rect 25044 2388 25096 2440
rect 47860 2456 47912 2508
rect 36728 2388 36780 2440
rect 48964 2388 49016 2440
rect 20260 2252 20312 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 662 49200 718 50000
rect 12898 49314 12954 50000
rect 12452 49286 12954 49314
rect 676 47122 704 49200
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 664 47116 716 47122
rect 664 47058 716 47064
rect 1584 47048 1636 47054
rect 1584 46990 1636 46996
rect 1596 24818 1624 46990
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 2410 38176 2466 38185
rect 2410 38111 2466 38120
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1492 24744 1544 24750
rect 1492 24686 1544 24692
rect 1504 2650 1532 24686
rect 2424 24682 2452 38111
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3424 25696 3476 25702
rect 3424 25638 3476 25644
rect 3436 25265 3464 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3422 25256 3478 25265
rect 3422 25191 3478 25200
rect 12452 24682 12480 49286
rect 12898 49200 12954 49286
rect 25134 49314 25190 50000
rect 25134 49286 25268 49314
rect 25134 49200 25190 49286
rect 25240 47054 25268 49286
rect 37370 49200 37426 50000
rect 49606 49200 49662 50000
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 25504 47184 25556 47190
rect 25504 47126 25556 47132
rect 25228 47048 25280 47054
rect 25228 46990 25280 46996
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 25044 37664 25096 37670
rect 25044 37606 25096 37612
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 25056 25906 25084 37606
rect 25044 25900 25096 25906
rect 25044 25842 25096 25848
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 25516 24818 25544 47126
rect 37384 46918 37412 49200
rect 37372 46912 37424 46918
rect 37372 46854 37424 46860
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 39316 25498 39344 46854
rect 49620 46102 49648 49200
rect 48136 46096 48188 46102
rect 48136 46038 48188 46044
rect 49608 46096 49660 46102
rect 49608 46038 49660 46044
rect 48044 37868 48096 37874
rect 48044 37810 48096 37816
rect 48056 37505 48084 37810
rect 48042 37496 48098 37505
rect 48042 37431 48098 37440
rect 48148 26234 48176 46038
rect 48056 26206 48176 26234
rect 39304 25492 39356 25498
rect 39304 25434 39356 25440
rect 41512 25288 41564 25294
rect 41512 25230 41564 25236
rect 41524 24886 41552 25230
rect 46756 25152 46808 25158
rect 46756 25094 46808 25100
rect 41512 24880 41564 24886
rect 41512 24822 41564 24828
rect 46768 24818 46796 25094
rect 25044 24812 25096 24818
rect 25044 24754 25096 24760
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 46756 24812 46808 24818
rect 46756 24754 46808 24760
rect 47860 24812 47912 24818
rect 47860 24754 47912 24760
rect 2412 24676 2464 24682
rect 2412 24618 2464 24624
rect 12440 24676 12492 24682
rect 12440 24618 12492 24624
rect 1768 24608 1820 24614
rect 1768 24550 1820 24556
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 1780 24206 1808 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 1768 24200 1820 24206
rect 1768 24142 1820 24148
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2792 12345 2820 24006
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 23492 16574 23520 24550
rect 23492 16546 24072 16574
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 2778 12336 2834 12345
rect 2778 12271 2834 12280
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 32 800 60 2382
rect 12268 800 12296 2382
rect 20272 2310 20300 7822
rect 20260 2304 20312 2310
rect 20260 2246 20312 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 18 0 74 800
rect 12254 0 12310 800
rect 24044 762 24072 16546
rect 25056 2446 25084 24754
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 47872 24410 47900 24754
rect 48056 24682 48084 26206
rect 48136 25288 48188 25294
rect 48136 25230 48188 25236
rect 48044 24676 48096 24682
rect 48044 24618 48096 24624
rect 48148 24585 48176 25230
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 47860 24404 47912 24410
rect 47860 24346 47912 24352
rect 47860 24200 47912 24206
rect 47860 24142 47912 24148
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 46386 11656 46442 11665
rect 46386 11591 46442 11600
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 46400 7750 46428 11591
rect 46388 7744 46440 7750
rect 46388 7686 46440 7692
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 47872 2514 47900 24142
rect 47860 2508 47912 2514
rect 47860 2450 47912 2456
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 48964 2440 49016 2446
rect 48964 2382 49016 2388
rect 24412 870 24532 898
rect 24412 762 24440 870
rect 24504 800 24532 870
rect 36740 800 36768 2382
rect 48976 800 49004 2382
rect 24044 734 24440 762
rect 24490 0 24546 800
rect 36726 0 36782 800
rect 48962 0 49018 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 2410 38120 2466 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 3422 25200 3478 25256
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 48042 37440 48098 37496
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 2778 12280 2834 12336
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 48134 24520 48190 24576
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 46386 11600 46442 11656
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
<< metal3 >>
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 0 38178 800 38208
rect 2405 38178 2471 38181
rect 0 38176 2471 38178
rect 0 38120 2410 38176
rect 2466 38120 2471 38176
rect 0 38118 2471 38120
rect 0 38088 800 38118
rect 2405 38115 2471 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 48037 37498 48103 37501
rect 49200 37498 50000 37528
rect 48037 37496 50000 37498
rect 48037 37440 48042 37496
rect 48098 37440 50000 37496
rect 48037 37438 50000 37440
rect 48037 37435 48103 37438
rect 49200 37408 50000 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25258 800 25288
rect 3417 25258 3483 25261
rect 0 25256 3483 25258
rect 0 25200 3422 25256
rect 3478 25200 3483 25256
rect 0 25198 3483 25200
rect 0 25168 800 25198
rect 3417 25195 3483 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 48129 24578 48195 24581
rect 49200 24578 50000 24608
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 49200 24488 50000 24518
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12338 800 12368
rect 2773 12338 2839 12341
rect 0 12336 2839 12338
rect 0 12280 2778 12336
rect 2834 12280 2839 12336
rect 0 12278 2839 12280
rect 0 12248 800 12278
rect 2773 12275 2839 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 46381 11658 46447 11661
rect 49200 11658 50000 11688
rect 46381 11656 50000 11658
rect 46381 11600 46386 11656
rect 46442 11600 50000 11656
rect 46381 11598 50000 11600
rect 46381 11595 46447 11598
rect 49200 11568 50000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_ef_sc_hd__decap_12  FILLER_0_6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1649977179
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1649977179
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1649977179
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1649977179
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1649977179
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1649977179
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1649977179
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1649977179
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1649977179
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1649977179
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1649977179
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1649977179
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1649977179
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_489
timestamp 1649977179
transform 1 0 46092 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1649977179
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_505
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_513
timestamp 1649977179
transform 1 0 48300 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1649977179
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1649977179
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1649977179
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1649977179
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1649977179
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1649977179
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1649977179
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1649977179
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1649977179
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1649977179
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1649977179
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1649977179
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_505
timestamp 1649977179
transform 1 0 47564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_513
timestamp 1649977179
transform 1 0 48300 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1649977179
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1649977179
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1649977179
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1649977179
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1649977179
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_513
timestamp 1649977179
transform 1 0 48300 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_513
timestamp 1649977179
transform 1 0 48300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_513
timestamp 1649977179
transform 1 0 48300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1649977179
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1649977179
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_513
timestamp 1649977179
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_257
timestamp 1649977179
transform 1 0 24748 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_262
timestamp 1649977179
transform 1 0 25208 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_274
timestamp 1649977179
transform 1 0 26312 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_286
timestamp 1649977179
transform 1 0 27416 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_298
timestamp 1649977179
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1649977179
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1649977179
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1649977179
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1649977179
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1649977179
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1649977179
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1649977179
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1649977179
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1649977179
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1649977179
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1649977179
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1649977179
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1649977179
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1649977179
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1649977179
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1649977179
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_513
timestamp 1649977179
transform 1 0 48300 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1649977179
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1649977179
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1649977179
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_513
timestamp 1649977179
transform 1 0 48300 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1649977179
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1649977179
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_513
timestamp 1649977179
transform 1 0 48300 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1649977179
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1649977179
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1649977179
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1649977179
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1649977179
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1649977179
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_513
timestamp 1649977179
transform 1 0 48300 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_513
timestamp 1649977179
transform 1 0 48300 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1649977179
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_513
timestamp 1649977179
transform 1 0 48300 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1649977179
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1649977179
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1649977179
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_513
timestamp 1649977179
transform 1 0 48300 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_513
timestamp 1649977179
transform 1 0 48300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_8
timestamp 1649977179
transform 1 0 1840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1649977179
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_507
timestamp 1649977179
transform 1 0 47748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1649977179
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_8
timestamp 1649977179
transform 1 0 1840 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_16
timestamp 1649977179
transform 1 0 2576 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_28
timestamp 1649977179
transform 1 0 3680 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_40
timestamp 1649977179
transform 1 0 4784 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1649977179
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1649977179
transform 1 0 25852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_277
timestamp 1649977179
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1649977179
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_437
timestamp 1649977179
transform 1 0 41308 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_443
timestamp 1649977179
transform 1 0 41860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_512
timestamp 1649977179
transform 1 0 48208 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_440
timestamp 1649977179
transform 1 0 41584 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_452
timestamp 1649977179
transform 1 0 42688 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_464
timestamp 1649977179
transform 1 0 43792 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1649977179
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_255
timestamp 1649977179
transform 1 0 24564 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_263
timestamp 1649977179
transform 1 0 25300 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1649977179
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_513
timestamp 1649977179
transform 1 0 48300 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1649977179
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1649977179
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1649977179
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1649977179
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1649977179
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1649977179
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1649977179
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1649977179
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_513
timestamp 1649977179
transform 1 0 48300 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1649977179
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1649977179
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1649977179
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1649977179
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1649977179
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1649977179
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1649977179
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1649977179
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1649977179
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1649977179
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1649977179
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1649977179
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1649977179
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1649977179
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1649977179
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1649977179
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1649977179
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1649977179
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1649977179
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_513
timestamp 1649977179
transform 1 0 48300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1649977179
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1649977179
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_513
timestamp 1649977179
transform 1 0 48300 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1649977179
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1649977179
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1649977179
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1649977179
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1649977179
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1649977179
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1649977179
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1649977179
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1649977179
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1649977179
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1649977179
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1649977179
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1649977179
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1649977179
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1649977179
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1649977179
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1649977179
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1649977179
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_512
timestamp 1649977179
transform 1 0 48208 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1649977179
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1649977179
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1649977179
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1649977179
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1649977179
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_513
timestamp 1649977179
transform 1 0 48300 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1649977179
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1649977179
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1649977179
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1649977179
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1649977179
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1649977179
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1649977179
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1649977179
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_513
timestamp 1649977179
transform 1 0 48300 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1649977179
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1649977179
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1649977179
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_513
timestamp 1649977179
transform 1 0 48300 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1649977179
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_513
timestamp 1649977179
transform 1 0 48300 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_513
timestamp 1649977179
transform 1 0 48300 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_513
timestamp 1649977179
transform 1 0 48300 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_513
timestamp 1649977179
transform 1 0 48300 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_513
timestamp 1649977179
transform 1 0 48300 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_13
timestamp 1649977179
transform 1 0 2300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_25
timestamp 1649977179
transform 1 0 3404 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_57
timestamp 1649977179
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_69
timestamp 1649977179
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1649977179
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_113
timestamp 1649977179
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_125
timestamp 1649977179
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1649977179
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_169
timestamp 1649977179
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_181
timestamp 1649977179
transform 1 0 17756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_193
timestamp 1649977179
transform 1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_225
timestamp 1649977179
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_237
timestamp 1649977179
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1649977179
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_261
timestamp 1649977179
transform 1 0 25116 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_281
timestamp 1649977179
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_293
timestamp 1649977179
transform 1 0 28060 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1649977179
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_337
timestamp 1649977179
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_349
timestamp 1649977179
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1649977179
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_393
timestamp 1649977179
transform 1 0 37260 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_405
timestamp 1649977179
transform 1 0 38364 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_417
timestamp 1649977179
transform 1 0 39468 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_449
timestamp 1649977179
transform 1 0 42412 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_461
timestamp 1649977179
transform 1 0 43516 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_473
timestamp 1649977179
transform 1 0 44620 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_505
timestamp 1649977179
transform 1 0 47564 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _00_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 47840 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _01_
timestamp 1649977179
transform -1 0 41860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _02_
timestamp 1649977179
transform -1 0 1840 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _03_
timestamp 1649977179
transform -1 0 25300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _04_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 41584 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1649977179
transform -1 0 1840 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1649977179
transform -1 0 24564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1649977179
transform 1 0 47840 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1649977179
transform 1 0 25484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1649977179
transform 1 0 2208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1649977179
transform -1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1649977179
transform 1 0 24840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 47932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 48208 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1649977179
transform -1 0 47104 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 25484 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 12604 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal3 s 49200 24488 50000 24608 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 662 49200 718 50000 0 FreeSans 224 90 0 0 io_in[1]
port 1 nsew signal input
flabel metal3 s 49200 37408 50000 37528 0 FreeSans 480 0 0 0 io_in[2]
port 2 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 io_in[3]
port 3 nsew signal input
flabel metal2 s 25134 49200 25190 50000 0 FreeSans 224 90 0 0 io_in[4]
port 4 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 io_in[5]
port 5 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 io_in[6]
port 6 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 io_in[7]
port 7 nsew signal input
flabel metal2 s 37370 49200 37426 50000 0 FreeSans 224 90 0 0 io_out[0]
port 8 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 io_out[1]
port 9 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 io_out[2]
port 10 nsew signal tristate
flabel metal2 s 49606 49200 49662 50000 0 FreeSans 224 90 0 0 io_out[3]
port 11 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 io_out[4]
port 12 nsew signal tristate
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 io_out[5]
port 13 nsew signal tristate
flabel metal2 s 12898 49200 12954 50000 0 FreeSans 224 90 0 0 io_out[6]
port 14 nsew signal tristate
flabel metal3 s 49200 11568 50000 11688 0 FreeSans 480 0 0 0 io_out[7]
port 15 nsew signal tristate
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
